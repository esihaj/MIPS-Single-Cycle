library verilog;
use verilog.vl_types.all;
entity test_stack is
end test_stack;
