library verilog;
use verilog.vl_types.all;
entity test_inst_memory is
end test_inst_memory;
