library verilog;
use verilog.vl_types.all;
entity test_data_memory is
end test_data_memory;
