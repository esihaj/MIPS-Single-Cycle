library verilog;
use verilog.vl_types.all;
entity test_reg_file is
end test_reg_file;
